module controlUnit # (
    parameter DATA_WIDTH = 32
)(
    input   logic       EQ,
    input   logic       instr,
    output  logic       RegWrite,
    output  logic       ALUctrl,
    output  logic       ALUsrc,
    output  logic       ImmSrc,
    output  logic       PCsrc
);


endmodule